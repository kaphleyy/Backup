//  verilog file

module start(a,b,c);
output c;
input a,b;

and G1(c,a,b);
endmodule;